`timescale 1ns / 1ps
`default_nettype none
//////////////////////////////////////////////////////////////////////////////////
// 
// Module Name:    encoder_to_rpm 
// Description: 
//
//////////////////////////////////////////////////////////////////////////////////
module encoder_to_rpm(cclk,rstb,a,b,rpm);
	//port definitions
	input  wire cclk;
	input  wire rstb;
	input  wire a;
	input  wire b;
	output wire [7:0] rpm;


endmodule
`default_nettype wire
